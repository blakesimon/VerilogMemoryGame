`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:42:21 12/02/2016 
// Design Name: 
// Module Name:    qini_count 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module qini_count(
    input qini,
    input qw,
    input qr,
    input clk,
    input reset,
    output flag
    );
	 reg count;
	 reg flag1;
always @(posedge clk)
begin
	
end

endmodule
