`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:29:21 12/01/2016 
// Design Name: 
// Module Name:    pb_scen 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module pb_scen(
    input yellow,
    input red,
    input blue,
    input green,
    output yel,
    output re,
    output blu,
    output gre,
    input reset,
    input clk
    );
always @(posedge clk)

endmodule
